module usb

interface ClassDriver {
	dev &Device
}
